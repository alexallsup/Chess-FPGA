// Btn Debouncer

module btn_debouncer(
	input CLK, input RESET,
	input Btn, output Btn_pulse);

endmodule