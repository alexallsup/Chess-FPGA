`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Alex Allsup & Kevin Wu
// 
// Create Date:    17:40:01 11/09/2016 
// Design Name: 
// Module Name:    game_logic 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module game_logic(
    input [255:0] board_input,
    output [5:0] board_out_addr,
    output [3:0] board_out_piece,
    input BtnL,
    input BtnU,
    input BtnR,
    input BtnD,
    input BtnC,
    output [5:0] highlight_square_addr
    );


endmodule
